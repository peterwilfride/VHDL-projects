--library ieee;
--use ieee.std_logic_1164.all;

--entity incrementer is
--	generic(b: in std_logic_vector(3 downto 0):="0001";
--				cin : in std_logic:="0");
--	port(a : in std_logic_vector(3 downto 0);
--			s : out std_logic_vector(3 downto 0);
--			cout : out std_logic);
--end incrementer;
--
--architecture behavior of incrementer is
--	component somador is
--	port(a, b, cin : in std_logic;
--		s, cout : out std_logic);
--	end component;
--	--signals
--	signal c: std_logic_vector(4 downto 0);
--	
--	begin
--		gen: for i in 0 to 3 generate
--			uut: somador port map (a(i), b(i), c(i), s(i), c(i+1));
--		end generate;
--		c(0) <= cin;
--		cout <= c(4);
--end behavior;