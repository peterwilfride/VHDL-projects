library verilog;
use verilog.vl_types.all;
entity wait_statement_vlg_sample_tst is
    port(
        clk_in          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end wait_statement_vlg_sample_tst;
