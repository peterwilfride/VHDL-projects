library verilog;
use verilog.vl_types.all;
entity comparator_4b_vlg_check_tst is
    port(
        aeqb            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end comparator_4b_vlg_check_tst;
