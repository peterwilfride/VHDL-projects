library verilog;
use verilog.vl_types.all;
entity wait_statement_vlg_check_tst is
    port(
        clk_out         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end wait_statement_vlg_check_tst;
