library ieee;
use ieee.std_logic_1164.all;

entity decrementer is
	generic(b: in std_logic_vector(3 downto 0):="0001";
				win : in std_logic:='0');
	port(a : in std_logic_vector(3 downto 0);
			s : out std_logic_vector(3 downto 0);
			wout : out std_logic);
end decrementer;

architecture behavior of decrementer is
	component subtrador_1b is
	port(a, b, win : in std_logic;
			s, wout : out std_logic);
	end component;
	--signals
	signal c: std_logic_vector(4 downto 0);
	
	begin
		gen: for i in 0 to 3 generate
			uut: subtrador_1b port map (a(i), b(i), c(i), s(i), c(i+1));
		end generate;
		c(0) <= win;
		wout <= c(4);
end behavior;