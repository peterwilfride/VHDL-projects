library verilog;
use verilog.vl_types.all;
entity wait_statement_vlg_vec_tst is
end wait_statement_vlg_vec_tst;
