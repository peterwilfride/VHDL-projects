entity display7seg is
port (s4, s3, s2, s1: in bit;
H7, H6, H5, H4, H3, H2, H1: out bit);
end display7seg;
architecture comportamento of display7seg is
begin
H1<=not(((not s4) and (not s3) and (not s2) and (not s1)) or ((not s4) and (not s3) and (s2) and (not s1)) or ((not s4) and (not s3) and (s2) and (s1)) or ((not s4) and (s3) and (not s2) and (s1)) or ((not s4) and (s3) and (s2) and (not s1)) or ((not s4) and (s3) and (s2) and (s1)) or ((s4) and (not s3) and (not s2) and (not s1)) or ((s4) and (not s3) and (not s2) and (s1)) or ((s4) and (not s3) and (s2) and (not s1)) or ((s4) and (s3) and (not s2) and (not s1)) or ((s4) and (s3) and (s2) and (not s1)) or ((s4) and (s3) and (s2) and (s1)));
H2<=not(((not s4) and (not s3) and (not s2) and (not s1))or  ((not s4) and (not s3) and (not s2) and (s1)) or ((not s4) and (not s3) and (s2) and (not s1)) or ((not s4) and (not s3) and (s2) and (s1)) or ((not s4) and (s3) and (not s2) and (not s1)) or ((not s4) and (s3) and (s2) and (s1)) or ((s4) and (not s3) and (not s2) and (not s1)) or ((s4) and (not s3) and (not s2) and (s1)) or ((s4) and (not s3) and (s2) and (not s1)) or ((s4) and (s3) and (not s2) and (s1)));
H3<=not (((not s4) and (not s3) and (not s2) and (not s1)) or ((not s4) and (not s3) and (not s2) and (s1)) or ((not s4) and (not s3) and (s2) and (s1)) or ((not s4) and (s3) and (not s2) and (not s1)) or ((not s4) and (s3) and (not s2) and (s1)) or ((not s4) and (s3) and (s2) and (not s1)) or ((not s4) and (s3) and (s2) and (s1)) or ((s4) and (not s3) and (not s2) and (not s1)) or ((s4) and (not s3) and (not s2) and (s1)) or ((s4) and (not s3) and (s2) and (not s1)) or ((s4) and (not s3) and (s2) and (s1)) or ((s4) and (s3) and (not s2) and (s1)));
H4<=not (((not s4) and (not s3) and (not s2) and (not s1)) or ((not s4) and (not s3) and (s2) and (not s1)) or ((not s4) and (not s3) and (s2) and (s1)) or ((not s4) and (s3) and (not s2) and (s1)) or ((not s4) and (s3) and (s2) and (not s1)) or ((s4) and (not s3) and (not s2) and (not s1)) or ((s4) and (not s3) and (not s2) and (s1)) or ((s4) and (not s3) and (s2) and (s1)) or ((s4) and (s3) and (not s2) and (not s1)) or ((s4) and (s3) and (not s2) and (s1)) or ((s4) and (s3) and (s2) and (not s1)));
H5<=not (((not s4) and (not s3) and (not s2) and (not s1)) or ((not s4) and (not s3) and (s2) and (not s1)) or ((not s4) and (s3) and (s2) and (not s1)) or ((s4) and (not s3) and (not s2) and (not s1)) or ((s4) and (not s3) and (s2) and (not s1)) or ((s4) and (not s3) and (s2) and (s1)) or ((s4) and (s3) and (not s2) and (not s1)) or ((s4) and (s3) and (not s2) and (s1)) or ((s4) and (s3) and (s2) and (not s1)) or ((s4) and (s3) and (s2) and (s1)));
H6<=not (((not s4) and (not s3) and (not s2) and (not s1)) or ((not s4) and (s3) and (not s2) and (not s1)) or ((not s4) and (s3) and (not s2) and (s1)) or ((not s4) and (s3) and (s2) and (not s1)) or ((s4) and (not s3) and (not s2) and (not s1)) or ((s4) and (not s3) and (not s2) and (s1)) or ((s4) and (not s3) and (s2) and (not s1)) or ((s4) and (not s3) and (s2) and (s1)) or ((s4) and (s3) and (not s2) and (not s1)) or ((s4) and (s3) and (s2) and (not s1)) or ((s4) and (s3) and (s2) and (s1)));
H7<=not (((not s4) and (not s3) and (s2) and (not s1)) or ((not s4) and (not s3) and (s2) and (s1)) or ((not s4) and (s3) and (not s2) and (not s1)) or ((not s4) and (s3) and (not s2) and (s1)) or ((not s4) and (s3) and (s2) and (not s1)) or ((s4) and (not s3) and (not s2) and (not s1)) or ((s4) and (not s3) and (not s2) and (s1)) or ((s4) and (not s3) and (s2) and (not s1)) or ((s4) and (not s3) and (s2) and (s1)) or ((s4) and (s3) and (not s2) and (s1)) or ((s4) and (s3) and (s2) and (not s1)) or ((s4) and (s3) and (s2) and (s1)));
end comportamento;