entity somador_quatro_bits is
	port(a: in bit_vector(3 downto 0);
	b: in bit_vector(3 downto 0);
	c0: in bit;
	s: out bit_vector(3 downto 0);
	c4: out bit);
end somador_quatro_bits;

architecture comportamento of somador_quatro_bits is

signal c3, c2, c1: bit;

begin
	s(0) <= a(0) xor b(0) xor c0;
	c1 <= ((a(0) xor b(0)) xor c0) or (a(0) and b(0));
	s(1) <= a(1) xor b(1) xor c0;
	c2 <= ((a(1) xor b(1)) xor c0) or (a(1) and b(1));
	s(2) <= a(2) xor b(2) xor c0;
	c3 <= ((a(2) xor b(2)) xor c0) or (a(2) and b(2));
	s(3) <= a(3) xor b(3) xor c0;
	c4 <= ((a(3) xor b(3)) xor c0) or (a(3) and b(3));
end comportamento;