library verilog;
use verilog.vl_types.all;
entity comparator_4b_vlg_vec_tst is
end comparator_4b_vlg_vec_tst;
