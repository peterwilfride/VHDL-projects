library verilog;
use verilog.vl_types.all;
entity timer_teste_vlg_vec_tst is
end timer_teste_vlg_vec_tst;
